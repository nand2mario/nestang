`ifndef _wishbone_slaves_vh_
`define _wishbone_slaves_vh_

parameter WISHBONE_SLAVE_ADDRESS_CHEATS_DATA  = 1

`endif