`define RES_720P
`define GW_IDE

package configPackage;  

    localparam SDRAM_DATA_WIDTH = 16;
    localparam SDRAM_ROW_WIDTH = 13;
    localparam SDRAM_COL_WIDTH = 9;
    localparam SDRAM_BANK_WIDTH = 2;

endpackage